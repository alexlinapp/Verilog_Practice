module addr_carry_param
    #(parameter N = 4)
    (
        input wire [N-1:0] a, b,
        output wire [N-1:0] sum,
        output wire cout
    );
    wire [N:0] sum_ext;
    assign sum_ext = {1'b0, a} + {1'b0, b};
    assign sum = sum_ext[N-1:0];
    assign cout = sum_ext[N];
endmodule
