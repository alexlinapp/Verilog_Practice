module top(
            input logic CLK_100MHZ, 
            input logic [3:0]

endmodule
