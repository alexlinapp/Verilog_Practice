class Transaction;








endclass : Transaction