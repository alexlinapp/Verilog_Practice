program automatic test();
    import abc::*;
    Transaction tr;
    // Test code
    initial begin
        $display("Program runs");
    end
    

endprogram


module top();
    test t1();
endmodule