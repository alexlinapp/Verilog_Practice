// Aysynchronous FIFO
//

module FIFO(

    );
endmodule
